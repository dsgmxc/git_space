module sine_wave #(
    parameter ACC_WIDTH = 32,		// 累加器宽度
    parameter ROM_WIDTH = 10,		// rom表深度
    parameter ANGLE_WIDTH = 16,		// 角度幅值位宽，q0.15格式
    parameter AMP_WIDTH = 16,		// 幅度比例位宽，q0.15格式
    parameter TIM_WIDTH = 16,		// 时间比例位宽 = 幅度比例位宽，q0.15格式
    parameter SEC_WIDTH = 3,		// 6个扇区
    parameter PHASE_WIDTH = 11		// 相位地址宽度 = rom表深度+1，数据对称点数翻倍
)(
    input  wire        clk,
    input  wire        rst_n,

    input  wire [ACC_WIDTH-1:0] phase_step,      // 相位步长，控制输出频率（Step = f*2^32/clk）
    input  wire signed [AMP_WIDTH-1:0] amplitude,         // 输出线电压的幅值 (Q15格式)(amplitude = A/V_DC*gen3)
	
    output reg [SEC_WIDTH-1:0] sectors,
    output reg [TIM_WIDTH-1:0] t1,
    output reg [TIM_WIDTH-1:0] t2,
    output reg  signed [AMP_WIDTH-1:0] va,       // A相电压 (Q15格式)
    output reg  signed [AMP_WIDTH-1:0] vb,       // B相电压 (Q15格式)
    output reg  signed [AMP_WIDTH-1:0] vc        // C相电压 (Q15格式)
);

    // --- 第1步：相位累加器 ---
    reg [ACC_WIDTH-1:0] phase_acc;      // 相位累加器

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            phase_acc <= 0;
        end else begin
            phase_acc <= phase_acc + phase_step;
        end
    end

    // --- 第2步：从ROM中查表获取三相余弦值 ---
    // 使用相位累加器的高位作为地址
wire [PHASE_WIDTH-1:0] rom_addr_a = phase_acc[ACC_WIDTH-1:ACC_WIDTH-PHASE_WIDTH];  
wire [PHASE_WIDTH-1:0] rom_addr_b = phase_acc[ACC_WIDTH-1:ACC_WIDTH-PHASE_WIDTH] + 11'd1365;  // 2^PHASE_WIDTH*2/3
wire [PHASE_WIDTH-1:0] rom_addr_c = phase_acc[ACC_WIDTH-1:ACC_WIDTH-PHASE_WIDTH] + 11'd682;  // 2^PHASE_WIDTH/3
wire over_a = rom_addr_a[PHASE_WIDTH-1] == 1'b1;  // 使用最高位判断
wire over_b = rom_addr_b[PHASE_WIDTH-1] == 1'b1;
wire over_c = rom_addr_c[PHASE_WIDTH-1] == 1'b1;
wire [PHASE_WIDTH - 2:0] addr_a = over_a ? ((1<<PHASE_WIDTH) - rom_addr_a[PHASE_WIDTH-1:0] - 1) : rom_addr_a[PHASE_WIDTH - 2:0];
wire [PHASE_WIDTH - 2:0] addr_b = over_b ? ((1<<PHASE_WIDTH) - rom_addr_b[PHASE_WIDTH-1:0] - 1) : rom_addr_b[PHASE_WIDTH - 2:0];
wire [PHASE_WIDTH - 2:0] addr_c = over_c ? ((1<<PHASE_WIDTH) - rom_addr_c[PHASE_WIDTH-1:0] - 1) : rom_addr_c[PHASE_WIDTH - 2:0];
reg signed [ANGLE_WIDTH-1:0] cos_table [0:(1<<ROM_WIDTH)-1];
initial begin
cos_table[0] = 16'sd32767;
cos_table[1] = 16'sd32767;
cos_table[2] = 16'sd32766;
cos_table[3] = 16'sd32766;
cos_table[4] = 16'sd32765;
cos_table[5] = 16'sd32763;
cos_table[6] = 16'sd32761;
cos_table[7] = 16'sd32759;
cos_table[8] = 16'sd32757;
cos_table[9] = 16'sd32754;
cos_table[10] = 16'sd32752;
cos_table[11] = 16'sd32748;
cos_table[12] = 16'sd32745;
cos_table[13] = 16'sd32741;
cos_table[14] = 16'sd32737;
cos_table[15] = 16'sd32732;
cos_table[16] = 16'sd32727;
cos_table[17] = 16'sd32722;
cos_table[18] = 16'sd32717;
cos_table[19] = 16'sd32711;
cos_table[20] = 16'sd32705;
cos_table[21] = 16'sd32699;
cos_table[22] = 16'sd32692;
cos_table[23] = 16'sd32685;
cos_table[24] = 16'sd32678;
cos_table[25] = 16'sd32670;
cos_table[26] = 16'sd32663;
cos_table[27] = 16'sd32654;
cos_table[28] = 16'sd32646;
cos_table[29] = 16'sd32637;
cos_table[30] = 16'sd32628;
cos_table[31] = 16'sd32619;
cos_table[32] = 16'sd32609;
cos_table[33] = 16'sd32599;
cos_table[34] = 16'sd32589;
cos_table[35] = 16'sd32578;
cos_table[36] = 16'sd32567;
cos_table[37] = 16'sd32556;
cos_table[38] = 16'sd32544;
cos_table[39] = 16'sd32532;
cos_table[40] = 16'sd32520;
cos_table[41] = 16'sd32508;
cos_table[42] = 16'sd32495;
cos_table[43] = 16'sd32482;
cos_table[44] = 16'sd32468;
cos_table[45] = 16'sd32455;
cos_table[46] = 16'sd32441;
cos_table[47] = 16'sd32426;
cos_table[48] = 16'sd32412;
cos_table[49] = 16'sd32397;
cos_table[50] = 16'sd32381;
cos_table[51] = 16'sd32366;
cos_table[52] = 16'sd32350;
cos_table[53] = 16'sd32334;
cos_table[54] = 16'sd32317;
cos_table[55] = 16'sd32301;
cos_table[56] = 16'sd32284;
cos_table[57] = 16'sd32266;
cos_table[58] = 16'sd32249;
cos_table[59] = 16'sd32231;
cos_table[60] = 16'sd32212;
cos_table[61] = 16'sd32194;
cos_table[62] = 16'sd32175;
cos_table[63] = 16'sd32156;
cos_table[64] = 16'sd32136;
cos_table[65] = 16'sd32116;
cos_table[66] = 16'sd32096;
cos_table[67] = 16'sd32076;
cos_table[68] = 16'sd32055;
cos_table[69] = 16'sd32034;
cos_table[70] = 16'sd32013;
cos_table[71] = 16'sd31991;
cos_table[72] = 16'sd31969;
cos_table[73] = 16'sd31947;
cos_table[74] = 16'sd31925;
cos_table[75] = 16'sd31902;
cos_table[76] = 16'sd31879;
cos_table[77] = 16'sd31855;
cos_table[78] = 16'sd31831;
cos_table[79] = 16'sd31807;
cos_table[80] = 16'sd31783;
cos_table[81] = 16'sd31758;
cos_table[82] = 16'sd31734;
cos_table[83] = 16'sd31708;
cos_table[84] = 16'sd31683;
cos_table[85] = 16'sd31657;
cos_table[86] = 16'sd31631;
cos_table[87] = 16'sd31604;
cos_table[88] = 16'sd31578;
cos_table[89] = 16'sd31551;
cos_table[90] = 16'sd31523;
cos_table[91] = 16'sd31496;
cos_table[92] = 16'sd31468;
cos_table[93] = 16'sd31440;
cos_table[94] = 16'sd31411;
cos_table[95] = 16'sd31382;
cos_table[96] = 16'sd31353;
cos_table[97] = 16'sd31324;
cos_table[98] = 16'sd31294;
cos_table[99] = 16'sd31264;
cos_table[100] = 16'sd31234;
cos_table[101] = 16'sd31203;
cos_table[102] = 16'sd31173;
cos_table[103] = 16'sd31141;
cos_table[104] = 16'sd31110;
cos_table[105] = 16'sd31078;
cos_table[106] = 16'sd31046;
cos_table[107] = 16'sd31014;
cos_table[108] = 16'sd30981;
cos_table[109] = 16'sd30948;
cos_table[110] = 16'sd30915;
cos_table[111] = 16'sd30882;
cos_table[112] = 16'sd30848;
cos_table[113] = 16'sd30814;
cos_table[114] = 16'sd30779;
cos_table[115] = 16'sd30745;
cos_table[116] = 16'sd30710;
cos_table[117] = 16'sd30675;
cos_table[118] = 16'sd30639;
cos_table[119] = 16'sd30603;
cos_table[120] = 16'sd30567;
cos_table[121] = 16'sd30531;
cos_table[122] = 16'sd30494;
cos_table[123] = 16'sd30457;
cos_table[124] = 16'sd30420;
cos_table[125] = 16'sd30382;
cos_table[126] = 16'sd30344;
cos_table[127] = 16'sd30306;
cos_table[128] = 16'sd30268;
cos_table[129] = 16'sd30229;
cos_table[130] = 16'sd30190;
cos_table[131] = 16'sd30151;
cos_table[132] = 16'sd30111;
cos_table[133] = 16'sd30072;
cos_table[134] = 16'sd30032;
cos_table[135] = 16'sd29991;
cos_table[136] = 16'sd29950;
cos_table[137] = 16'sd29910;
cos_table[138] = 16'sd29868;
cos_table[139] = 16'sd29827;
cos_table[140] = 16'sd29785;
cos_table[141] = 16'sd29743;
cos_table[142] = 16'sd29701;
cos_table[143] = 16'sd29658;
cos_table[144] = 16'sd29615;
cos_table[145] = 16'sd29572;
cos_table[146] = 16'sd29528;
cos_table[147] = 16'sd29485;
cos_table[148] = 16'sd29440;
cos_table[149] = 16'sd29396;
cos_table[150] = 16'sd29352;
cos_table[151] = 16'sd29307;
cos_table[152] = 16'sd29262;
cos_table[153] = 16'sd29216;
cos_table[154] = 16'sd29170;
cos_table[155] = 16'sd29124;
cos_table[156] = 16'sd29078;
cos_table[157] = 16'sd29032;
cos_table[158] = 16'sd28985;
cos_table[159] = 16'sd28938;
cos_table[160] = 16'sd28890;
cos_table[161] = 16'sd28843;
cos_table[162] = 16'sd28795;
cos_table[163] = 16'sd28747;
cos_table[164] = 16'sd28698;
cos_table[165] = 16'sd28650;
cos_table[166] = 16'sd28601;
cos_table[167] = 16'sd28552;
cos_table[168] = 16'sd28502;
cos_table[169] = 16'sd28452;
cos_table[170] = 16'sd28402;
cos_table[171] = 16'sd28352;
cos_table[172] = 16'sd28301;
cos_table[173] = 16'sd28250;
cos_table[174] = 16'sd28199;
cos_table[175] = 16'sd28148;
cos_table[176] = 16'sd28096;
cos_table[177] = 16'sd28044;
cos_table[178] = 16'sd27992;
cos_table[179] = 16'sd27940;
cos_table[180] = 16'sd27887;
cos_table[181] = 16'sd27834;
cos_table[182] = 16'sd27781;
cos_table[183] = 16'sd27727;
cos_table[184] = 16'sd27674;
cos_table[185] = 16'sd27620;
cos_table[186] = 16'sd27565;
cos_table[187] = 16'sd27511;
cos_table[188] = 16'sd27456;
cos_table[189] = 16'sd27401;
cos_table[190] = 16'sd27346;
cos_table[191] = 16'sd27290;
cos_table[192] = 16'sd27234;
cos_table[193] = 16'sd27178;
cos_table[194] = 16'sd27122;
cos_table[195] = 16'sd27065;
cos_table[196] = 16'sd27008;
cos_table[197] = 16'sd26951;
cos_table[198] = 16'sd26894;
cos_table[199] = 16'sd26836;
cos_table[200] = 16'sd26778;
cos_table[201] = 16'sd26720;
cos_table[202] = 16'sd26662;
cos_table[203] = 16'sd26603;
cos_table[204] = 16'sd26545;
cos_table[205] = 16'sd26485;
cos_table[206] = 16'sd26426;
cos_table[207] = 16'sd26366;
cos_table[208] = 16'sd26307;
cos_table[209] = 16'sd26246;
cos_table[210] = 16'sd26186;
cos_table[211] = 16'sd26125;
cos_table[212] = 16'sd26065;
cos_table[213] = 16'sd26003;
cos_table[214] = 16'sd25942;
cos_table[215] = 16'sd25881;
cos_table[216] = 16'sd25819;
cos_table[217] = 16'sd25757;
cos_table[218] = 16'sd25694;
cos_table[219] = 16'sd25632;
cos_table[220] = 16'sd25569;
cos_table[221] = 16'sd25506;
cos_table[222] = 16'sd25443;
cos_table[223] = 16'sd25379;
cos_table[224] = 16'sd25315;
cos_table[225] = 16'sd25251;
cos_table[226] = 16'sd25187;
cos_table[227] = 16'sd25123;
cos_table[228] = 16'sd25058;
cos_table[229] = 16'sd24993;
cos_table[230] = 16'sd24928;
cos_table[231] = 16'sd24862;
cos_table[232] = 16'sd24797;
cos_table[233] = 16'sd24731;
cos_table[234] = 16'sd24665;
cos_table[235] = 16'sd24598;
cos_table[236] = 16'sd24532;
cos_table[237] = 16'sd24465;
cos_table[238] = 16'sd24398;
cos_table[239] = 16'sd24330;
cos_table[240] = 16'sd24263;
cos_table[241] = 16'sd24195;
cos_table[242] = 16'sd24127;
cos_table[243] = 16'sd24059;
cos_table[244] = 16'sd23991;
cos_table[245] = 16'sd23922;
cos_table[246] = 16'sd23853;
cos_table[247] = 16'sd23784;
cos_table[248] = 16'sd23715;
cos_table[249] = 16'sd23645;
cos_table[250] = 16'sd23575;
cos_table[251] = 16'sd23505;
cos_table[252] = 16'sd23435;
cos_table[253] = 16'sd23365;
cos_table[254] = 16'sd23294;
cos_table[255] = 16'sd23223;
cos_table[256] = 16'sd23152;
cos_table[257] = 16'sd23081;
cos_table[258] = 16'sd23009;
cos_table[259] = 16'sd22937;
cos_table[260] = 16'sd22865;
cos_table[261] = 16'sd22793;
cos_table[262] = 16'sd22721;
cos_table[263] = 16'sd22648;
cos_table[264] = 16'sd22575;
cos_table[265] = 16'sd22502;
cos_table[266] = 16'sd22429;
cos_table[267] = 16'sd22356;
cos_table[268] = 16'sd22282;
cos_table[269] = 16'sd22208;
cos_table[270] = 16'sd22134;
cos_table[271] = 16'sd22060;
cos_table[272] = 16'sd21985;
cos_table[273] = 16'sd21910;
cos_table[274] = 16'sd21836;
cos_table[275] = 16'sd21760;
cos_table[276] = 16'sd21685;
cos_table[277] = 16'sd21610;
cos_table[278] = 16'sd21534;
cos_table[279] = 16'sd21458;
cos_table[280] = 16'sd21382;
cos_table[281] = 16'sd21305;
cos_table[282] = 16'sd21229;
cos_table[283] = 16'sd21152;
cos_table[284] = 16'sd21075;
cos_table[285] = 16'sd20998;
cos_table[286] = 16'sd20921;
cos_table[287] = 16'sd20843;
cos_table[288] = 16'sd20765;
cos_table[289] = 16'sd20687;
cos_table[290] = 16'sd20609;
cos_table[291] = 16'sd20531;
cos_table[292] = 16'sd20452;
cos_table[293] = 16'sd20374;
cos_table[294] = 16'sd20295;
cos_table[295] = 16'sd20216;
cos_table[296] = 16'sd20136;
cos_table[297] = 16'sd20057;
cos_table[298] = 16'sd19977;
cos_table[299] = 16'sd19897;
cos_table[300] = 16'sd19817;
cos_table[301] = 16'sd19737;
cos_table[302] = 16'sd19657;
cos_table[303] = 16'sd19576;
cos_table[304] = 16'sd19495;
cos_table[305] = 16'sd19414;
cos_table[306] = 16'sd19333;
cos_table[307] = 16'sd19252;
cos_table[308] = 16'sd19170;
cos_table[309] = 16'sd19089;
cos_table[310] = 16'sd19007;
cos_table[311] = 16'sd18925;
cos_table[312] = 16'sd18842;
cos_table[313] = 16'sd18760;
cos_table[314] = 16'sd18677;
cos_table[315] = 16'sd18595;
cos_table[316] = 16'sd18512;
cos_table[317] = 16'sd18429;
cos_table[318] = 16'sd18345;
cos_table[319] = 16'sd18262;
cos_table[320] = 16'sd18178;
cos_table[321] = 16'sd18094;
cos_table[322] = 16'sd18010;
cos_table[323] = 16'sd17926;
cos_table[324] = 16'sd17842;
cos_table[325] = 16'sd17757;
cos_table[326] = 16'sd17673;
cos_table[327] = 16'sd17588;
cos_table[328] = 16'sd17503;
cos_table[329] = 16'sd17418;
cos_table[330] = 16'sd17333;
cos_table[331] = 16'sd17247;
cos_table[332] = 16'sd17161;
cos_table[333] = 16'sd17076;
cos_table[334] = 16'sd16990;
cos_table[335] = 16'sd16904;
cos_table[336] = 16'sd16817;
cos_table[337] = 16'sd16731;
cos_table[338] = 16'sd16644;
cos_table[339] = 16'sd16557;
cos_table[340] = 16'sd16471;
cos_table[341] = 16'sd16384;
cos_table[342] = 16'sd16296;
cos_table[343] = 16'sd16209;
cos_table[344] = 16'sd16121;
cos_table[345] = 16'sd16034;
cos_table[346] = 16'sd15946;
cos_table[347] = 16'sd15858;
cos_table[348] = 16'sd15770;
cos_table[349] = 16'sd15681;
cos_table[350] = 16'sd15593;
cos_table[351] = 16'sd15504;
cos_table[352] = 16'sd15416;
cos_table[353] = 16'sd15327;
cos_table[354] = 16'sd15238;
cos_table[355] = 16'sd15149;
cos_table[356] = 16'sd15059;
cos_table[357] = 16'sd14970;
cos_table[358] = 16'sd14880;
cos_table[359] = 16'sd14791;
cos_table[360] = 16'sd14701;
cos_table[361] = 16'sd14611;
cos_table[362] = 16'sd14521;
cos_table[363] = 16'sd14430;
cos_table[364] = 16'sd14340;
cos_table[365] = 16'sd14249;
cos_table[366] = 16'sd14159;
cos_table[367] = 16'sd14068;
cos_table[368] = 16'sd13977;
cos_table[369] = 16'sd13886;
cos_table[370] = 16'sd13795;
cos_table[371] = 16'sd13703;
cos_table[372] = 16'sd13612;
cos_table[373] = 16'sd13520;
cos_table[374] = 16'sd13429;
cos_table[375] = 16'sd13337;
cos_table[376] = 16'sd13245;
cos_table[377] = 16'sd13153;
cos_table[378] = 16'sd13060;
cos_table[379] = 16'sd12968;
cos_table[380] = 16'sd12876;
cos_table[381] = 16'sd12783;
cos_table[382] = 16'sd12690;
cos_table[383] = 16'sd12597;
cos_table[384] = 16'sd12505;
cos_table[385] = 16'sd12411;
cos_table[386] = 16'sd12318;
cos_table[387] = 16'sd12225;
cos_table[388] = 16'sd12132;
cos_table[389] = 16'sd12038;
cos_table[390] = 16'sd11944;
cos_table[391] = 16'sd11851;
cos_table[392] = 16'sd11757;
cos_table[393] = 16'sd11663;
cos_table[394] = 16'sd11569;
cos_table[395] = 16'sd11474;
cos_table[396] = 16'sd11380;
cos_table[397] = 16'sd11286;
cos_table[398] = 16'sd11191;
cos_table[399] = 16'sd11097;
cos_table[400] = 16'sd11002;
cos_table[401] = 16'sd10907;
cos_table[402] = 16'sd10812;
cos_table[403] = 16'sd10717;
cos_table[404] = 16'sd10622;
cos_table[405] = 16'sd10527;
cos_table[406] = 16'sd10431;
cos_table[407] = 16'sd10336;
cos_table[408] = 16'sd10240;
cos_table[409] = 16'sd10145;
cos_table[410] = 16'sd10049;
cos_table[411] = 16'sd9953;
cos_table[412] = 16'sd9857;
cos_table[413] = 16'sd9761;
cos_table[414] = 16'sd9665;
cos_table[415] = 16'sd9569;
cos_table[416] = 16'sd9473;
cos_table[417] = 16'sd9376;
cos_table[418] = 16'sd9280;
cos_table[419] = 16'sd9183;
cos_table[420] = 16'sd9087;
cos_table[421] = 16'sd8990;
cos_table[422] = 16'sd8893;
cos_table[423] = 16'sd8796;
cos_table[424] = 16'sd8699;
cos_table[425] = 16'sd8602;
cos_table[426] = 16'sd8505;
cos_table[427] = 16'sd8408;
cos_table[428] = 16'sd8311;
cos_table[429] = 16'sd8213;
cos_table[430] = 16'sd8116;
cos_table[431] = 16'sd8018;
cos_table[432] = 16'sd7921;
cos_table[433] = 16'sd7823;
cos_table[434] = 16'sd7725;
cos_table[435] = 16'sd7627;
cos_table[436] = 16'sd7529;
cos_table[437] = 16'sd7431;
cos_table[438] = 16'sd7333;
cos_table[439] = 16'sd7235;
cos_table[440] = 16'sd7137;
cos_table[441] = 16'sd7039;
cos_table[442] = 16'sd6941;
cos_table[443] = 16'sd6842;
cos_table[444] = 16'sd6744;
cos_table[445] = 16'sd6645;
cos_table[446] = 16'sd6547;
cos_table[447] = 16'sd6448;
cos_table[448] = 16'sd6349;
cos_table[449] = 16'sd6251;
cos_table[450] = 16'sd6152;
cos_table[451] = 16'sd6053;
cos_table[452] = 16'sd5954;
cos_table[453] = 16'sd5855;
cos_table[454] = 16'sd5756;
cos_table[455] = 16'sd5657;
cos_table[456] = 16'sd5558;
cos_table[457] = 16'sd5459;
cos_table[458] = 16'sd5359;
cos_table[459] = 16'sd5260;
cos_table[460] = 16'sd5161;
cos_table[461] = 16'sd5061;
cos_table[462] = 16'sd4962;
cos_table[463] = 16'sd4862;
cos_table[464] = 16'sd4763;
cos_table[465] = 16'sd4663;
cos_table[466] = 16'sd4564;
cos_table[467] = 16'sd4464;
cos_table[468] = 16'sd4364;
cos_table[469] = 16'sd4264;
cos_table[470] = 16'sd4165;
cos_table[471] = 16'sd4065;
cos_table[472] = 16'sd3965;
cos_table[473] = 16'sd3865;
cos_table[474] = 16'sd3765;
cos_table[475] = 16'sd3665;
cos_table[476] = 16'sd3565;
cos_table[477] = 16'sd3465;
cos_table[478] = 16'sd3365;
cos_table[479] = 16'sd3265;
cos_table[480] = 16'sd3165;
cos_table[481] = 16'sd3065;
cos_table[482] = 16'sd2964;
cos_table[483] = 16'sd2864;
cos_table[484] = 16'sd2764;
cos_table[485] = 16'sd2664;
cos_table[486] = 16'sd2563;
cos_table[487] = 16'sd2463;
cos_table[488] = 16'sd2363;
cos_table[489] = 16'sd2262;
cos_table[490] = 16'sd2162;
cos_table[491] = 16'sd2061;
cos_table[492] = 16'sd1961;
cos_table[493] = 16'sd1861;
cos_table[494] = 16'sd1760;
cos_table[495] = 16'sd1660;
cos_table[496] = 16'sd1559;
cos_table[497] = 16'sd1459;
cos_table[498] = 16'sd1358;
cos_table[499] = 16'sd1258;
cos_table[500] = 16'sd1157;
cos_table[501] = 16'sd1056;
cos_table[502] = 16'sd956;
cos_table[503] = 16'sd855;
cos_table[504] = 16'sd755;
cos_table[505] = 16'sd654;
cos_table[506] = 16'sd553;
cos_table[507] = 16'sd453;
cos_table[508] = 16'sd352;
cos_table[509] = 16'sd252;
cos_table[510] = 16'sd151;
cos_table[511] = 16'sd50;
cos_table[512] = -16'sd50;
cos_table[513] = -16'sd151;
    cos_table[514] = -16'sd252;
    cos_table[515] = -16'sd352;
    cos_table[516] = -16'sd453;
    cos_table[517] = -16'sd553;
    cos_table[518] = -16'sd654;
    cos_table[519] = -16'sd755;
    cos_table[520] = -16'sd855;
    cos_table[521] = -16'sd956;
    cos_table[522] = -16'sd1056;
    cos_table[523] = -16'sd1157;
    cos_table[524] = -16'sd1258;
    cos_table[525] = -16'sd1358;
    cos_table[526] = -16'sd1459;
    cos_table[527] = -16'sd1559;
    cos_table[528] = -16'sd1660;
    cos_table[529] = -16'sd1760;
    cos_table[530] = -16'sd1861;
    cos_table[531] = -16'sd1961;
    cos_table[532] = -16'sd2061;
    cos_table[533] = -16'sd2162;
    cos_table[534] = -16'sd2262;
    cos_table[535] = -16'sd2363;
    cos_table[536] = -16'sd2463;
    cos_table[537] = -16'sd2563;
    cos_table[538] = -16'sd2664;
    cos_table[539] = -16'sd2764;
    cos_table[540] = -16'sd2864;
    cos_table[541] = -16'sd2964;
    cos_table[542] = -16'sd3065;
    cos_table[543] = -16'sd3165;
    cos_table[544] = -16'sd3265;
    cos_table[545] = -16'sd3365;
    cos_table[546] = -16'sd3465;
    cos_table[547] = -16'sd3565;
    cos_table[548] = -16'sd3665;
    cos_table[549] = -16'sd3765;
    cos_table[550] = -16'sd3865;
    cos_table[551] = -16'sd3965;
    cos_table[552] = -16'sd4065;
    cos_table[553] = -16'sd4165;
    cos_table[554] = -16'sd4264;
    cos_table[555] = -16'sd4364;
    cos_table[556] = -16'sd4464;
    cos_table[557] = -16'sd4564;
    cos_table[558] = -16'sd4663;
    cos_table[559] = -16'sd4763;
    cos_table[560] = -16'sd4862;
    cos_table[561] = -16'sd4962;
    cos_table[562] = -16'sd5061;
    cos_table[563] = -16'sd5161;
    cos_table[564] = -16'sd5260;
    cos_table[565] = -16'sd5359;
    cos_table[566] = -16'sd5459;
    cos_table[567] = -16'sd5558;
    cos_table[568] = -16'sd5657;
    cos_table[569] = -16'sd5756;
    cos_table[570] = -16'sd5855;
    cos_table[571] = -16'sd5954;
    cos_table[572] = -16'sd6053;
    cos_table[573] = -16'sd6152;
    cos_table[574] = -16'sd6251;
    cos_table[575] = -16'sd6349;
    cos_table[576] = -16'sd6448;
    cos_table[577] = -16'sd6547;
    cos_table[578] = -16'sd6645;
    cos_table[579] = -16'sd6744;
    cos_table[580] = -16'sd6842;
    cos_table[581] = -16'sd6941;
    cos_table[582] = -16'sd7039;
    cos_table[583] = -16'sd7137;
    cos_table[584] = -16'sd7235;
    cos_table[585] = -16'sd7333;
    cos_table[586] = -16'sd7431;
    cos_table[587] = -16'sd7529;
    cos_table[588] = -16'sd7627;
    cos_table[589] = -16'sd7725;
    cos_table[590] = -16'sd7823;
    cos_table[591] = -16'sd7921;
    cos_table[592] = -16'sd8018;
    cos_table[593] = -16'sd8116;
    cos_table[594] = -16'sd8213;
    cos_table[595] = -16'sd8311;
    cos_table[596] = -16'sd8408;
    cos_table[597] = -16'sd8505;
    cos_table[598] = -16'sd8602;
    cos_table[599] = -16'sd8699;
    cos_table[600] = -16'sd8796;
    cos_table[601] = -16'sd8893;
    cos_table[602] = -16'sd8990;
    cos_table[603] = -16'sd9087;
    cos_table[604] = -16'sd9183;
    cos_table[605] = -16'sd9280;
    cos_table[606] = -16'sd9376;
    cos_table[607] = -16'sd9473;
    cos_table[608] = -16'sd9569;
    cos_table[609] = -16'sd9665;
    cos_table[610] = -16'sd9761;
    cos_table[611] = -16'sd9857;
    cos_table[612] = -16'sd9953;
    cos_table[613] = -16'sd10049;
    cos_table[614] = -16'sd10145;
    cos_table[615] = -16'sd10240;
    cos_table[616] = -16'sd10336;
    cos_table[617] = -16'sd10431;
    cos_table[618] = -16'sd10527;
    cos_table[619] = -16'sd10622;
    cos_table[620] = -16'sd10717;
    cos_table[621] = -16'sd10812;
    cos_table[622] = -16'sd10907;
    cos_table[623] = -16'sd11002;
    cos_table[624] = -16'sd11097;
    cos_table[625] = -16'sd11191;
    cos_table[626] = -16'sd11286;
    cos_table[627] = -16'sd11380;
    cos_table[628] = -16'sd11474;
    cos_table[629] = -16'sd11569;
    cos_table[630] = -16'sd11663;
    cos_table[631] = -16'sd11757;
    cos_table[632] = -16'sd11851;
    cos_table[633] = -16'sd11944;
    cos_table[634] = -16'sd12038;
    cos_table[635] = -16'sd12132;
    cos_table[636] = -16'sd12225;
    cos_table[637] = -16'sd12318;
    cos_table[638] = -16'sd12411;
    cos_table[639] = -16'sd12505;
    cos_table[640] = -16'sd12597;
    cos_table[641] = -16'sd12690;
    cos_table[642] = -16'sd12783;
    cos_table[643] = -16'sd12876;
    cos_table[644] = -16'sd12968;
    cos_table[645] = -16'sd13060;
    cos_table[646] = -16'sd13153;
    cos_table[647] = -16'sd13245;
    cos_table[648] = -16'sd13337;
    cos_table[649] = -16'sd13429;
    cos_table[650] = -16'sd13520;
    cos_table[651] = -16'sd13612;
    cos_table[652] = -16'sd13703;
    cos_table[653] = -16'sd13795;
    cos_table[654] = -16'sd13886;
    cos_table[655] = -16'sd13977;
    cos_table[656] = -16'sd14068;
    cos_table[657] = -16'sd14159;
    cos_table[658] = -16'sd14249;
    cos_table[659] = -16'sd14340;
    cos_table[660] = -16'sd14430;
    cos_table[661] = -16'sd14521;
    cos_table[662] = -16'sd14611;
    cos_table[663] = -16'sd14701;
    cos_table[664] = -16'sd14791;
    cos_table[665] = -16'sd14880;
    cos_table[666] = -16'sd14970;
    cos_table[667] = -16'sd15059;
    cos_table[668] = -16'sd15149;
    cos_table[669] = -16'sd15238;
    cos_table[670] = -16'sd15327;
    cos_table[671] = -16'sd15416;
    cos_table[672] = -16'sd15504;
    cos_table[673] = -16'sd15593;
    cos_table[674] = -16'sd15681;
    cos_table[675] = -16'sd15770;
    cos_table[676] = -16'sd15858;
    cos_table[677] = -16'sd15946;
    cos_table[678] = -16'sd16034;
    cos_table[679] = -16'sd16121;
    cos_table[680] = -16'sd16209;
    cos_table[681] = -16'sd16296;
    cos_table[682] = -16'sd16383;
    cos_table[683] = -16'sd16471;
    cos_table[684] = -16'sd16557;
    cos_table[685] = -16'sd16644;
    cos_table[686] = -16'sd16731;
    cos_table[687] = -16'sd16817;
    cos_table[688] = -16'sd16904;
    cos_table[689] = -16'sd16990;
    cos_table[690] = -16'sd17076;
    cos_table[691] = -16'sd17161;
    cos_table[692] = -16'sd17247;
    cos_table[693] = -16'sd17333;
    cos_table[694] = -16'sd17418;
    cos_table[695] = -16'sd17503;
    cos_table[696] = -16'sd17588;
    cos_table[697] = -16'sd17673;
    cos_table[698] = -16'sd17757;
    cos_table[699] = -16'sd17842;
    cos_table[700] = -16'sd17926;
    cos_table[701] = -16'sd18010;
    cos_table[702] = -16'sd18094;
    cos_table[703] = -16'sd18178;
    cos_table[704] = -16'sd18262;
    cos_table[705] = -16'sd18345;
    cos_table[706] = -16'sd18429;
    cos_table[707] = -16'sd18512;
    cos_table[708] = -16'sd18595;
    cos_table[709] = -16'sd18677;
    cos_table[710] = -16'sd18760;
    cos_table[711] = -16'sd18842;
    cos_table[712] = -16'sd18925;
    cos_table[713] = -16'sd19007;
    cos_table[714] = -16'sd19089;
    cos_table[715] = -16'sd19170;
    cos_table[716] = -16'sd19252;
    cos_table[717] = -16'sd19333;
    cos_table[718] = -16'sd19414;
    cos_table[719] = -16'sd19495;
    cos_table[720] = -16'sd19576;
    cos_table[721] = -16'sd19657;
    cos_table[722] = -16'sd19737;
    cos_table[723] = -16'sd19817;
    cos_table[724] = -16'sd19897;
    cos_table[725] = -16'sd19977;
    cos_table[726] = -16'sd20057;
    cos_table[727] = -16'sd20136;
    cos_table[728] = -16'sd20216;
    cos_table[729] = -16'sd20295;
    cos_table[730] = -16'sd20374;
    cos_table[731] = -16'sd20452;
    cos_table[732] = -16'sd20531;
    cos_table[733] = -16'sd20609;
    cos_table[734] = -16'sd20687;
    cos_table[735] = -16'sd20765;
    cos_table[736] = -16'sd20843;
    cos_table[737] = -16'sd20921;
    cos_table[738] = -16'sd20998;
    cos_table[739] = -16'sd21075;
    cos_table[740] = -16'sd21152;
    cos_table[741] = -16'sd21229;
    cos_table[742] = -16'sd21305;
    cos_table[743] = -16'sd21382;
    cos_table[744] = -16'sd21458;
    cos_table[745] = -16'sd21534;
    cos_table[746] = -16'sd21610;
    cos_table[747] = -16'sd21685;
    cos_table[748] = -16'sd21760;
    cos_table[749] = -16'sd21836;
    cos_table[750] = -16'sd21910;
    cos_table[751] = -16'sd21985;
    cos_table[752] = -16'sd22060;
    cos_table[753] = -16'sd22134;
    cos_table[754] = -16'sd22208;
    cos_table[755] = -16'sd22282;
    cos_table[756] = -16'sd22356;
    cos_table[757] = -16'sd22429;
    cos_table[758] = -16'sd22502;
    cos_table[759] = -16'sd22575;
    cos_table[760] = -16'sd22648;
    cos_table[761] = -16'sd22721;
    cos_table[762] = -16'sd22793;
    cos_table[763] = -16'sd22865;
    cos_table[764] = -16'sd22937;
    cos_table[765] = -16'sd23009;
    cos_table[766] = -16'sd23081;
    cos_table[767] = -16'sd23152;
    cos_table[768] = -16'sd23223;
    cos_table[769] = -16'sd23294;
    cos_table[770] = -16'sd23365;
    cos_table[771] = -16'sd23435;
    cos_table[772] = -16'sd23505;
    cos_table[773] = -16'sd23575;
    cos_table[774] = -16'sd23645;
    cos_table[775] = -16'sd23715;
    cos_table[776] = -16'sd23784;
    cos_table[777] = -16'sd23853;
    cos_table[778] = -16'sd23922;
    cos_table[779] = -16'sd23991;
    cos_table[780] = -16'sd24059;
    cos_table[781] = -16'sd24127;
    cos_table[782] = -16'sd24195;
    cos_table[783] = -16'sd24263;
    cos_table[784] = -16'sd24330;
    cos_table[785] = -16'sd24398;
    cos_table[786] = -16'sd24465;
    cos_table[787] = -16'sd24532;
    cos_table[788] = -16'sd24598;
    cos_table[789] = -16'sd24665;
    cos_table[790] = -16'sd24731;
    cos_table[791] = -16'sd24797;
    cos_table[792] = -16'sd24862;
    cos_table[793] = -16'sd24928;
    cos_table[794] = -16'sd24993;
    cos_table[795] = -16'sd25058;
    cos_table[796] = -16'sd25123;
    cos_table[797] = -16'sd25187;
    cos_table[798] = -16'sd25251;
    cos_table[799] = -16'sd25315;
    cos_table[800] = -16'sd25379;
    cos_table[801] = -16'sd25443;
    cos_table[802] = -16'sd25506;
    cos_table[803] = -16'sd25569;
    cos_table[804] = -16'sd25632;
    cos_table[805] = -16'sd25694;
    cos_table[806] = -16'sd25757;
    cos_table[807] = -16'sd25819;
    cos_table[808] = -16'sd25881;
    cos_table[809] = -16'sd25942;
    cos_table[810] = -16'sd26003;
    cos_table[811] = -16'sd26065;
    cos_table[812] = -16'sd26125;
    cos_table[813] = -16'sd26186;
    cos_table[814] = -16'sd26246;
    cos_table[815] = -16'sd26307;
    cos_table[816] = -16'sd26366;
    cos_table[817] = -16'sd26426;
    cos_table[818] = -16'sd26485;
    cos_table[819] = -16'sd26545;
    cos_table[820] = -16'sd26603;
    cos_table[821] = -16'sd26662;
    cos_table[822] = -16'sd26720;
    cos_table[823] = -16'sd26778;
    cos_table[824] = -16'sd26836;
    cos_table[825] = -16'sd26894;
    cos_table[826] = -16'sd26951;
    cos_table[827] = -16'sd27008;
    cos_table[828] = -16'sd27065;
    cos_table[829] = -16'sd27122;
    cos_table[830] = -16'sd27178;
    cos_table[831] = -16'sd27234;
    cos_table[832] = -16'sd27290;
    cos_table[833] = -16'sd27346;
    cos_table[834] = -16'sd27401;
    cos_table[835] = -16'sd27456;
    cos_table[836] = -16'sd27511;
    cos_table[837] = -16'sd27565;
    cos_table[838] = -16'sd27620;
    cos_table[839] = -16'sd27674;
    cos_table[840] = -16'sd27727;
    cos_table[841] = -16'sd27781;
    cos_table[842] = -16'sd27834;
    cos_table[843] = -16'sd27887;
    cos_table[844] = -16'sd27940;
    cos_table[845] = -16'sd27992;
    cos_table[846] = -16'sd28044;
    cos_table[847] = -16'sd28096;
    cos_table[848] = -16'sd28148;
    cos_table[849] = -16'sd28199;
    cos_table[850] = -16'sd28250;
    cos_table[851] = -16'sd28301;
    cos_table[852] = -16'sd28352;
    cos_table[853] = -16'sd28402;
    cos_table[854] = -16'sd28452;
    cos_table[855] = -16'sd28502;
    cos_table[856] = -16'sd28552;
    cos_table[857] = -16'sd28601;
    cos_table[858] = -16'sd28650;
    cos_table[859] = -16'sd28698;
    cos_table[860] = -16'sd28747;
    cos_table[861] = -16'sd28795;
    cos_table[862] = -16'sd28843;
    cos_table[863] = -16'sd28890;
    cos_table[864] = -16'sd28938;
    cos_table[865] = -16'sd28985;
    cos_table[866] = -16'sd29032;
    cos_table[867] = -16'sd29078;
    cos_table[868] = -16'sd29124;
    cos_table[869] = -16'sd29170;
    cos_table[870] = -16'sd29216;
    cos_table[871] = -16'sd29262;
    cos_table[872] = -16'sd29307;
    cos_table[873] = -16'sd29352;
    cos_table[874] = -16'sd29396;
    cos_table[875] = -16'sd29440;
    cos_table[876] = -16'sd29485;
    cos_table[877] = -16'sd29528;
    cos_table[878] = -16'sd29572;
    cos_table[879] = -16'sd29615;
    cos_table[880] = -16'sd29658;
    cos_table[881] = -16'sd29701;
    cos_table[882] = -16'sd29743;
    cos_table[883] = -16'sd29785;
    cos_table[884] = -16'sd29827;
    cos_table[885] = -16'sd29868;
    cos_table[886] = -16'sd29910;
    cos_table[887] = -16'sd29950;
    cos_table[888] = -16'sd29991;
    cos_table[889] = -16'sd30032;
    cos_table[890] = -16'sd30072;
    cos_table[891] = -16'sd30111;
    cos_table[892] = -16'sd30151;
    cos_table[893] = -16'sd30190;
    cos_table[894] = -16'sd30229;
    cos_table[895] = -16'sd30268;
    cos_table[896] = -16'sd30306;
    cos_table[897] = -16'sd30344;
    cos_table[898] = -16'sd30382;
    cos_table[899] = -16'sd30420;
    cos_table[900] = -16'sd30457;
    cos_table[901] = -16'sd30494;
    cos_table[902] = -16'sd30531;
    cos_table[903] = -16'sd30567;
    cos_table[904] = -16'sd30603;
    cos_table[905] = -16'sd30639;
    cos_table[906] = -16'sd30675;
    cos_table[907] = -16'sd30710;
    cos_table[908] = -16'sd30745;
    cos_table[909] = -16'sd30779;
    cos_table[910] = -16'sd30814;
    cos_table[911] = -16'sd30848;
    cos_table[912] = -16'sd30882;
    cos_table[913] = -16'sd30915;
    cos_table[914] = -16'sd30948;
    cos_table[915] = -16'sd30981;
    cos_table[916] = -16'sd31014;
    cos_table[917] = -16'sd31046;
    cos_table[918] = -16'sd31078;
    cos_table[919] = -16'sd31110;
    cos_table[920] = -16'sd31141;
    cos_table[921] = -16'sd31173;
    cos_table[922] = -16'sd31203;
    cos_table[923] = -16'sd31234;
    cos_table[924] = -16'sd31264;
    cos_table[925] = -16'sd31294;
    cos_table[926] = -16'sd31324;
    cos_table[927] = -16'sd31353;
    cos_table[928] = -16'sd31382;
    cos_table[929] = -16'sd31411;
    cos_table[930] = -16'sd31440;
    cos_table[931] = -16'sd31468;
    cos_table[932] = -16'sd31496;
    cos_table[933] = -16'sd31523;
    cos_table[934] = -16'sd31551;
    cos_table[935] = -16'sd31578;
    cos_table[936] = -16'sd31604;
    cos_table[937] = -16'sd31631;
    cos_table[938] = -16'sd31657;
    cos_table[939] = -16'sd31683;
    cos_table[940] = -16'sd31708;
    cos_table[941] = -16'sd31734;
    cos_table[942] = -16'sd31758;
    cos_table[943] = -16'sd31783;
    cos_table[944] = -16'sd31807;
    cos_table[945] = -16'sd31831;
    cos_table[946] = -16'sd31855;
    cos_table[947] = -16'sd31879;
    cos_table[948] = -16'sd31902;
    cos_table[949] = -16'sd31925;
    cos_table[950] = -16'sd31947;
    cos_table[951] = -16'sd31969;
    cos_table[952] = -16'sd31991;
    cos_table[953] = -16'sd32013;
    cos_table[954] = -16'sd32034;
    cos_table[955] = -16'sd32055;
    cos_table[956] = -16'sd32076;
    cos_table[957] = -16'sd32096;
    cos_table[958] = -16'sd32116;
    cos_table[959] = -16'sd32136;
    cos_table[960] = -16'sd32156;
    cos_table[961] = -16'sd32175;
    cos_table[962] = -16'sd32194;
    cos_table[963] = -16'sd32212;
    cos_table[964] = -16'sd32231;
    cos_table[965] = -16'sd32249;
    cos_table[966] = -16'sd32266;
    cos_table[967] = -16'sd32284;
    cos_table[968] = -16'sd32301;
    cos_table[969] = -16'sd32317;
    cos_table[970] = -16'sd32334;
    cos_table[971] = -16'sd32350;
    cos_table[972] = -16'sd32366;
    cos_table[973] = -16'sd32381;
    cos_table[974] = -16'sd32397;
    cos_table[975] = -16'sd32412;
    cos_table[976] = -16'sd32426;
    cos_table[977] = -16'sd32441;
    cos_table[978] = -16'sd32455;
    cos_table[979] = -16'sd32468;
    cos_table[980] = -16'sd32482;
    cos_table[981] = -16'sd32495;
    cos_table[982] = -16'sd32508;
    cos_table[983] = -16'sd32520;
    cos_table[984] = -16'sd32532;
    cos_table[985] = -16'sd32544;
    cos_table[986] = -16'sd32556;
    cos_table[987] = -16'sd32567;
    cos_table[988] = -16'sd32578;
    cos_table[989] = -16'sd32589;
    cos_table[990] = -16'sd32599;
    cos_table[991] = -16'sd32609;
    cos_table[992] = -16'sd32619;
    cos_table[993] = -16'sd32628;
    cos_table[994] = -16'sd32637;
    cos_table[995] = -16'sd32646;
    cos_table[996] = -16'sd32654;
    cos_table[997] = -16'sd32663;
    cos_table[998] = -16'sd32670;
    cos_table[999] = -16'sd32678;
    cos_table[1000] = -16'sd32685;
    cos_table[1001] = -16'sd32692;
    cos_table[1002] = -16'sd32699;
    cos_table[1003] = -16'sd32705;
    cos_table[1004] = -16'sd32711;
    cos_table[1005] = -16'sd32717;
    cos_table[1006] = -16'sd32722;
    cos_table[1007] = -16'sd32727;
    cos_table[1008] = -16'sd32732;
    cos_table[1009] = -16'sd32737;
    cos_table[1010] = -16'sd32741;
    cos_table[1011] = -16'sd32745;
    cos_table[1012] = -16'sd32748;
    cos_table[1013] = -16'sd32752;
    cos_table[1014] = -16'sd32754;
    cos_table[1015] = -16'sd32757;
    cos_table[1016] = -16'sd32759;
    cos_table[1017] = -16'sd32761;
    cos_table[1018] = -16'sd32763;
    cos_table[1019] = -16'sd32765;
    cos_table[1020] = -16'sd32766;
    cos_table[1021] = -16'sd32766;
    cos_table[1022] = -16'sd32767;
    cos_table[1023] = -16'sd32767;
end
    wire signed [ANGLE_WIDTH + AMP_WIDTH - 1:0] cos_val_a = cos_table[addr_a] * amplitude;
    wire signed [ANGLE_WIDTH + AMP_WIDTH - 1:0] cos_val_b = cos_table[addr_b] * amplitude;
    wire signed [ANGLE_WIDTH + AMP_WIDTH - 1:0] cos_val_c = cos_table[addr_c] * amplitude;
    reg [PHASE_WIDTH - 1:0] phase;
    // --- 第3步：乘以幅值，得到最终输出 ---
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            va <= 0;
            vb <= 0;
            vc <= 0;
            phase <= 0;
        end else begin
            va <= cos_val_a[ANGLE_WIDTH+AMP_WIDTH-2:ANGLE_WIDTH-1];
            vb <= cos_val_b[ANGLE_WIDTH+AMP_WIDTH-2:ANGLE_WIDTH-1];
            vc <= cos_val_c[ANGLE_WIDTH+AMP_WIDTH-2:ANGLE_WIDTH-1];
            phase <= rom_addr_a;
        end
    end
    
    // --- 第4步：扇区判断 ---
    // 临时变量用于组合逻辑计算
    wire signed [AMP_WIDTH - 1:0] v_ab = va - vb;
    wire signed [AMP_WIDTH - 1:0] v_bc = vb - vc;
    wire signed [AMP_WIDTH - 1:0] v_ca = vc - va; 
    reg signed [TIM_WIDTH - 1:0] t1_temp, t2_temp;
    reg [SEC_WIDTH-1:0] sectors_temp;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            t1 <= 0;
            t2 <= 0;
            sectors <= 1;
            t1_temp <= 0;
            t2_temp <= 0;
            sectors_temp <= 1;
        end else begin
            // 根据相位判断扇区（使用新的512点边界）
            if (phase < 11'd344) begin          // 扇区1: 0°-60°
                sectors_temp <= 3'd1;
                t1_temp = v_ab;  
                t2_temp = v_bc;
            end 
            else if (phase < 11'd684) begin     // 扇区2: 60°-120°
                sectors_temp <= 3'd2;
                t1_temp = -v_ca;
                t2_temp = -v_ab;
            end 
            else if (phase < 11'd1024) begin    // 扇区3: 120°-180°
                sectors_temp <= 3'd3;
                t1_temp = v_bc;
                t2_temp = v_ca;
            end 
            else if (phase < 11'd1364) begin    // 扇区4: 180°-240°
                sectors_temp <= 3'd4;
                t1_temp = -v_ab;
                t2_temp = -v_bc;
            end 
            else if (phase < 11'd1704) begin    // 扇区5: 240°-300°
                sectors_temp <= 3'd5;
                t1_temp = v_ca;
                t2_temp = v_ab;
            end 
            else begin                        // 扇区6: 300°-360°
                sectors_temp <= 3'd6;
                t1_temp = -v_bc;
                t2_temp = -v_ca;
            end
            // 负值限制为0
            t1 <= (t1_temp[TIM_WIDTH - 1]) ? 0 : t1_temp;
            t2 <= (t2_temp[TIM_WIDTH - 1]) ? 0 : t2_temp;
            sectors <= sectors_temp;
        end
    end

endmodule



